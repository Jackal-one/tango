module top (
    input i_clk,
    input i_rstn
);
    
endmodule